module demo

