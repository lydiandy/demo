module controller

import demo
import model

pub fn create_product(c demo.Context) {

}