module middleware

pub fn gzip() Middleware {
}
