module middleware

pub fn request_id() Middleware {
}
