// after create table,insert the init data
module main

fn main() {
}
