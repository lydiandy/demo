module middleware

pub fn timeout() Middleware {
}
