module demo

pub struct Router {
}
