module middleware

pub fn session() Middleware {
}
