module middleware

pub fn recover() {
}
