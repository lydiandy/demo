module demo

type Middleware fn(*Context)

type Handler fn(*Context)

// type Middleware fn(Handler) Handler 




