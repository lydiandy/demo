module middleware

pub fn compress() Middleware {
}
