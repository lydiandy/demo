module model

pub struct Product {
}
