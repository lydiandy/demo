module mobile

import demo

pub fn login(c demo.Context) {
}
