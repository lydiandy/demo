module middleware

pub fn recover() Middleware {
}
