module middleware

pub fn body_limit() Middleware {
}
