module middleware

pub fn static_file() Middleware {
}
