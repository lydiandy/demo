module middleware

pub fn static_file(path string) {
	
}