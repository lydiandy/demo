module middleware

pub fn cors() Middleware {
}
