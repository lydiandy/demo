module test

pub fn test_app() {
	
}