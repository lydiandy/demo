module middleware

pub fn redirect() Middleware {
}
