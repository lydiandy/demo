module controller

import demo
import model

pub fn get_user_list(c demo.Context) {
}

pub fn get_user_detail(c demo.Context) {
}

pub fn create_user(c demo.Context) {
}

pub fn edit_user(c demo.Context) {
}

pub fn remove_user(c demo.Context) {
}
