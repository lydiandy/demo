module middleware

pub fn logger() Middleware {
}
