module model

module model

pub struct User {
	
}