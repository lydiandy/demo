module logger

//usage:
//import demo.logger
//app.use(logger.new(cfg))

pub struct Config() {

}

pub fn new(cfg Config) {
	
}


