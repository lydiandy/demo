module middleware

pub fn favicon() Middleware {
}
