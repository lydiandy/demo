module middleware

pub fn jwt() Middleware {
}
